.title KiCad schematic
.include "models/BZX84C4V7.spice.txt"
.include "models/C2012C0G2A102J060AA_p.mod"
.include "models/CGJ4C2C0G2A101J060AA_p.mod"
.include "models/FMMT597.spice.txt"
.include "models/SMAZ15.spice.txt"
.include "models/ZXCT1010.spice.txt"
XU4 0 /COCM /PWR_IN /SN ZXCT1010
XU5 /PWR_IN /SN CGJ4C2C0G2A101J060AA_p
R5 /SN /PWR_OUT 10k
R6 /PWR_IN /PWR_OUT 0.04
XU3 /BASE /PWR_IN SMAZ15
Q1 /COLLECTOR /BASE /COCM FMMT597
R3 0 /BASE 1.5Meg
R1 /OUT /COLLECTOR 100
R2 /COLLECTOR 0 4.99k
XU2 /OUT 0 C2012C0G2A102J060AA_p
XU1 0 /OUT DI_BZX84C4V7
I1 /PWR_OUT 0 {ILOAD}
V1 /PWR_IN 0 {VSOURCE}
R7 /PWR_IN /PWR_OUT 0.04
R4 /COLLECTOR 0 4.99k
.end
